module mycpu_top(
    input  wire        aresetn,
    input  wire        aclk,

    output wire [3 :0] arid,
    output wire [31:0] araddr, 
    output wire [7 :0] arlen,  
    output wire [2 :0] arsize, 
    output wire [1 :0] arburst,
    output wire [1 :0] arlock, 
    output wire [3 :0] arcache,
    output wire [2 :0] arprot, 
    output wire        arvalid,
    input  wire        arready,
    input  wire [3 :0] rid,    
    input  wire [31:0] rdata,  
    input  wire [1 :0] rresp,  
    input  wire        rlast,  
    input  wire        rvalid, 
    output wire        rready, 
    output wire [3 :0] awid,   
    output wire [31:0] awaddr, 
    output wire [7 :0] awlen,  
    output wire [2 :0] awsize, 
    output wire [1 :0] awburst,
    output wire [1 :0] awlock, 
    output wire [3 :0] awcache,
    output wire [2 :0] awprot, 
    output wire        awvalid,
    input  wire        awready,
    output wire [3 :0] wid,    
    output wire [31:0] wdata,  
    output wire [3 :0] wstrb,  
    output wire        wlast,  
    output wire        wvalid, 
    input  wire        wready, 
    input  wire [3 :0] bid,    
    input  wire [1 :0] bresp,  
    input  wire        bvalid, 
    output wire        bready, 

    output wire [31:0] debug_wb_pc,
    output wire [ 3:0] debug_wb_rf_wen,
    output wire [ 4:0] debug_wb_rf_wnum,
    output wire [31:0] debug_wb_rf_wdata

);
widsnoy_cpu mycpu(
    .clock                      (aclk),
    .reset                      (~aresetn),
    .io_axi_arid                (arid),
    .io_axi_araddr              (araddr),
    .io_axi_arlen               (arlen),
    .io_axi_arsize              (arsize),
    .io_axi_arburst             (arburst),
    .io_axi_arlock              (arlock),
    .io_axi_arcache             (arcache),
    .io_axi_arprot              (arprot),
    .io_axi_arvalid             (arvalid),
    .io_axi_arready             (arready),
    .io_axi_rid                 (rid),
    .io_axi_rready              (rready),
    .io_axi_rdata               (rdata),
    .io_axi_rvalid              (rvalid),
    .io_axi_awid                (awid),
    .io_axi_awaddr              (awaddr),
    .io_axi_awlen               (awlen),
    .io_axi_awsize              (awsize),
    .io_axi_awburst             (awburst),
    .io_axi_awlock              (awlock),
    .io_axi_awcache             (awcache),
    .io_axi_awprot              (awprot),
    .io_axi_awvalid             (awvalid),
    .io_axi_awready             (awready),
    .io_axi_wid                 (wid),
    .io_axi_wdata               (wdata),
    .io_axi_wstrb               (wstrb),
    .io_axi_wlast               (wlast),
    .io_axi_wvalid              (wvalid),
    .io_axi_wready              (wready),
    .io_axi_bvalid              (bvalid),
    .io_axi_bready              (bready),
    .io_debug_wb_pc             (debug_wb_pc),
    .io_debug_wb_rf_wen         (debug_wb_rf_wen),    
    .io_debug_wb_rf_wnum        (debug_wb_rf_wnum),        
    .io_debug_wb_rf_wdata       (debug_wb_rf_wdata)       
);
endmodule