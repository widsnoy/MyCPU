module mycpu_top(

);
widsnoy_cpu mycpu(

);
endmodule